module uurisc #(
    parameters
) (
    port_list
);
    
endmodule